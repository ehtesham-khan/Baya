module top
(input wire gclk, gresetn, pclk, presetn, clk_phase,
			cpu_clk, cpu_resetn, dmx_clk, dmx_resetn);

endmodule

