module master ( bus_intf.master intf_master, input clock ); 
endmodule
