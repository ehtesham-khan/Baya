module slave ( bus_intf.slave intf_slave, input clock, output out1 ); 
endmodule
