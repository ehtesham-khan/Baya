module dmxwrp (
				input wire rst_n,dmx_clk,gresetn,gclk,presetn,pclk,clk_phase,
				input wire ts_clk_a,fr_ts_sync_a,fr_ts_dvalid_a,
				input wire [7:0] fr_ts_di_a,
				input wire fr_ts_derr_a,
				apb_bus apb_dmx			,
				axi_bus.axi_master_aw axi_dmx	,
				output wire out_int
);
dmx			u_dmx					(
				.rst_n					(rst_n					),
				.dmx_clk				(dmx_clk				),
				.gresetn				(gresetn				),
				.gclk					(gclk					),
				.presetn				(presetn				),
				.pclk					(pclk					),
				.clk_phase				(clk_phase				),
				.ts_clk_a				(ts_clk_a				),
				.fr_ts_sync_a			(fr_ts_sync_a			),
				.fr_ts_dvalid_a			(fr_ts_dvalid_a			),
				.fr_ts_di_a				(fr_ts_di_a				),
				.fr_ts_derr_a			(fr_ts_derr_a			),
				.penable				(apb_dmx.penable		),
				.psel					(apb_dmx.psel			),
				.pwrite					(apb_dmx.pwrite			),
				.paddr					(apb_dmx.paddr[13:2]	),
				.pwdata					(apb_dmx.pwdata			),
				.prdata					(apb_dmx.prdata			),
				.pready					(apb_dmx.pready			),
				.aid_dmx				(axi_dmx.aid			),
				.axi_addr_dmx			(axi_dmx.aaddr			),
				.avalid_dmx				(axi_dmx.avalid			),
				.awrite_dmx				(axi_dmx.awrite			),
				.alen_dmx				(axi_dmx.alen			),
				.asize_dmx				(axi_dmx.asize			),
				.aburst_dmx				(axi_dmx.aburst			),
				.wid_dmx				(axi_dmx.wid			),
				.wdata_dmx				(axi_dmx.wdata			),
				.wstrb_dmx				(axi_dmx.wstrb			),
				.wlast_dmx				(axi_dmx.wlast			),
				.wvalid_dmx				(axi_dmx.wvalid			),
				.aready_dmx				(axi_dmx.aready			),
				.wready_dmx				(axi_dmx.wready			),
				.out_int				(out_int				) 
);
endmodule
