-- ****************************************************************************
-- ** Description: types.vhd
-- ** Author:      The SPIRIT Consortium
-- ** 
-- ** 
-- ** Revision:    $Revision: 1.1 $
-- ** Date:        $Date: 2014/12/27 22:48:30 $
-- ** 
-- ** Copyright (c) 2008, 2009 The SPIRIT Consortium.
-- ** 
-- ** This work forms part of a deliverable of The SPIRIT Consortium.
-- ** 
-- ** Use of these materials are governed by the legal terms and conditions
-- ** outlined in the disclaimer available from www.spiritconsortium.org.
-- ** 
-- ** This source file is provided on an AS IS basis.  The SPIRIT
-- ** Consortium disclaims any warranty express or implied including
-- ** any warranty of merchantability and fitness for use for a
-- ** particular purpose.
-- ** 
-- ** The user of the source file shall indemnify and hold The SPIRIT
-- ** Consortium and its members harmless from any damages or liability.
-- ** Users are requested to provide feedback to The SPIRIT Consortium
-- ** using either mailto:feedback@lists.spiritconsortium.org or the forms at 
-- ** http://www.spiritconsortium.org/about/contact_us/
-- ** 
-- ** This file may be copied, and distributed, with or without
-- ** modifications; this notice must be included on any copy.
-- ****************************************************************************

-----------------------------------------------------------------------------
-- Entity:      types
-- File:        types.vhd
-- Author:      SPIRIT IP-XACT
-- Description: Package with type declarations 
------------------------------------------------------------------------------
  
library IEEE;
use IEEE.std_logic_1164.all;

package types is


subtype clk_type is std_logic;
subtype dac_word_type is std_logic_vector(23 downto 0);


end;

