module MySoC( clk, out1 );
	input clk;
	output out1;
endmodule 
