module B(
        a,
        b,
        c
    );
    output[7:0] a;
    output[7:0] b;
    input[7:0] c;
endmodule 
