module C(
        a,
        b,
        c
    );
    input[7:0] a;
    output[7:0] b;
    output[7:0] c;
endmodule 
