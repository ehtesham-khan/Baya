module buswrp(
	input wire gclk, gresetn,cpu_clk,cpu_resetn,clk_phase,
	axi_bus.axi_slave_ar axi_audio,
	axi_bus.axi_slave_aw axi_demux,
	axi_bus.axi_slave axi_gdma,
	axi_bus.axi_master axi_ddr,
	apb_bus.apb_master1 apb_m,
	apb_bus.apb_master2 apb_s0,
	apb_bus.apb_master2 apb_s1,
	output wire sram_cen,
	output wire [7:0] sram_wen,
	output wire [9:0] sram_addr,
	output wire [63:0] sram_datain,
	input wire [63:0] sram_dataout
);

bus u_bus(
        .gclk					(gclk				),
        .gresetn				(gresetn			),
        .cpu_clk				(cpu_clk			),
        .cpu_resetn				(cpu_resetn			),
        .clk_phase				(clk_phase			),
        .aid_audioout			(axi_audio.aid		),
        .axi_addr_audioout		(axi_audio.aaddr	),
        .avalid_audioout		(axi_audio.avalid	),
        .awrite_audioout		(axi_audio.awrite	),
        .alen_audioout			(axi_audio.alen		),
        .asize_audioout			(axi_audio.asize	),
        .aburst_audioout		(axi_audio.aburst	),
        .rready_audioout		(axi_audio.rready	),
        .aready_audioout		(axi_audio.aready	),
        .rid_audioout			(axi_audio.rid		),
        .rdata_audioout			(axi_audio.rdata	),
        .rlast_audioout			(axi_audio.rlast	),
        .rvalid_audioout		(axi_audio.rvalid	),
        .aid_gdma				(axi_gdma.aid		),
        .axi_addr_gdma			(axi_gdma.aaddr		),
        .avalid_gdma			(axi_gdma.avalid	),
        .awrite_gdma			(axi_gdma.awrite	),
        .alen_gdma				(axi_gdma.alen		),
        .asize_gdma				(axi_gdma.asize		),
        .aburst_gdma			(axi_gdma.aburst	),
        .wid_gdma				(axi_gdma.wid		),
        .wdata_gdma				(axi_gdma.wdata		),
        .wstrb_gdma				(axi_gdma.wstrb		),
        .wlast_gdma				(axi_gdma.wlast		),
        .wvalid_gdma			(axi_gdma.wvalid	),
        .rready_gdma			(axi_gdma.rready	),
        .aready_gdma			(axi_gdma.aready	),
        .wready_gdma			(axi_gdma.wready	),
        .rid_gdma				(axi_gdma.rid		),
        .rdata_gdma				(axi_gdma.rdata		),
        .rlast_gdma				(axi_gdma.rlast		),
        .rvalid_gdma			(axi_gdma.rvalid	),
        .aid_demux				(axi_demux.aid		),
        .axi_addr_demux			(axi_demux.aaddr	),
        .avalid_demux			(axi_demux.avalid	),
        .awrite_demux			(axi_demux.awrite	),
        .alen_demux				(axi_demux.alen		),
        .asize_demux			(axi_demux.asize	),
        .aburst_demux			(axi_demux.aburst	),
        .wid_demux				(axi_demux.wid		),
        .wdata_demux			(axi_demux.wdata	),
        .wstrb_demux			(axi_demux.wstrb	),
        .wlast_demux			(axi_demux.wlast	),
        .wvalid_demux			(axi_demux.wvalid	),
        .aready_demux			(axi_demux.aready	),
        .wready_demux			(axi_demux.wready	),
        .aid_ddr				(axi_ddr.aid		),
        .axi_addr_ddr			(axi_ddr.aaddr		),
        .avalid_ddr				(axi_ddr.avalid		),
        .awrite_ddr				(axi_ddr.awrite		),
        .alen_ddr				(axi_ddr.alen		),
        .aburst_ddr				(axi_ddr.aburst		),
        .wid_ddr				(axi_ddr.wid		),
        .wdata_ddr				(axi_ddr.wdata		),
        .wstrb_ddr				(axi_ddr.wstrb		),
        .wlast_ddr				(axi_ddr.wlast		),
        .wvalid_ddr				(axi_ddr.wvalid		),
        .rready_ddr				(axi_ddr.rready		),
        .aready_ddr				(axi_ddr.aready		),
        .wready_ddr				(axi_ddr.wready		),
        .rid_ddr				(axi_ddr.rid		),
        .rdata_ddr				(axi_ddr.rdata		),
        .rlast_ddr				(axi_ddr.rlast		),
        .rvalid_ddr				(axi_ddr.rvalid		),
        .paddr					(apb_m.paddr		),
        .penable				(apb_m.penable		),
        .pwrite					(apb_m.pwrite		),
        .pwdata					(apb_m.pwdata		),
        .psel0					(apb_s0.psel		),
        .psel1					(apb_s1.psel		),
        .pready0				(apb_s0.pready		),
        .pready1				(apb_s1.pready		),
        .prdata0				(apb_s0.prdata		),
        .prdata1				(apb_s1.prdata		),
		.sram_cen				(sram_cen			),
		.sram_wen				(sram_wen			),
		.sram_addr				(sram_addr			),
		.sram_datain			(sram_datain		),
		.sram_dataout			(sram_dataout		)
);
endmodule
